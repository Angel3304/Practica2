library ieee; 
use ieee.std_logic_1164.all; 
use ieee.std_logic_arith.all; 
use ieee.std_logic_unsigned.all; ------------------------------------------------------------------------------------------------ 
entity Procesador_Top is 
 port( 
  clk : in std_logic; 
  switch : in std_logic_vector(1 downto 0); 
  Displays : out std_logic_vector(3 downto 0); 
  Segmentos : out std_logic_vector(7 downto 0) 
 ); 
end entity; 
------------------------------------------------------------------------------------------------- 
architecture behavioral of Procesador_Top is 
 
 --Señales 
 signal pc_aux : std_logic_vector(5 downto 0); 
 signal flag_loop : std_logic := '0'; 
 signal flag_start1 : std_logic := '0'; 
 signal flag_start2 : std_logic := '0'; 
 signal flag_start3 : std_logic := '0'; 
  
 signal rom_output_aux : std_logic_vector(21 downto 0); 
  
 signal output_ex_aux : std_logic_vector(9 downto 0); 
 signal flag_zero_aux : std_logic; 
 signal flag_signo_aux : std_logic; 
 signal flag_acarreo_aux : std_logic; 
 signal flag_overflow_aux : std_logic; 
  
 signal output_bcd_aux : std_logic_vector(15 downto 0); 
  
 signal output_uni_aux : std_logic_vector(7 downto 0); 
 signal output_dec_aux : std_logic_vector(7 downto 0); 
 signal output_cen_aux : std_logic_vector(7 downto 0); 
 signal output_mil_aux : std_logic_vector(7 downto 0); 
  
 signal cuenta : integer range 0 to 100000; 
 signal Seleccion : std_logic_vector(1 downto 0) := "00"; 
 signal Mostrar : std_logic_vector(3 downto 0) := "0000"; 
 ------------------------------------------------- 
  
 --Declaracion de omponentes 
  --Componente Rom 
 component Memoria_Instrucciones 
  port( 
   input : in std_logic_vector(5 downto 0); 
   output : out std_logic_vector(21 downto 0) 
 ); 
 end component; 
  
  --Componente Execute 
 component Unidad_Ejecucion 
  port( 
  input_ex : in std_logic_vector(21 downto 0); 
  output_ex : out std_logic_vector(9 downto 0); 
  flag_zero : out std_logic; 
  flag_signo : out std_logic; 
  flag_acarreo : out std_logic; 
  flag_overflow : out std_logic 
 ); 
 end component; 
 
 --Componente BCD 
 component Converti 
  Port ( 
   S : in  std_logic_vector(11 downto 0); 
   output_bcd : out std_logic_vector(15 downto 0) 
  ); 
 end component; 
 
 --Componente Mux display del resultado 
 component Parte2 
  Port(    
   input : in std_logic_vector(3 downto 0); 
   output: out std_logic_vector(7 downto 0) 
  ); 
 end component; -------------------------------------------------------------------------------------- 
begin 
 
 process(clk) 
 begin 
  case switch is 
   when "00" => 
    if flag_start1 = '0' then  
     if flag_loop = '0' then  
      pc_aux <= "000000"; 
      flag_loop <= '1'; 
     else 
      pc_aux <= pc_aux + '1'; 
     end if; 
    end if; 
   when "01" =>  
    if flag_start2 = '0' then  
     if flag_loop = '0' then  
      pc_aux <= "001010"; 
      flag_loop <= '1'; 
     else 
      pc_aux <= pc_aux + '1'; 
     end if; 
    end if; 
   when "10" =>  
    if flag_start3 = '0' then  
     if flag_loop = '0' then  
      pc_aux <= "010110"; 
      flag_loop <= '1'; 
     else 
      pc_aux <= pc_aux + '1'; 
     end if; 
    end if; 
   when "11" => 
    pc_aux <= "111111"; 
  end case; 
 end process; 
       
 process(clk) 
 begin 
  if rising_edge(clk) then  
   if pc_aux = "001001" then  
    flag_start1 <= '1'; 
    flag_start2 <= '0'; 
    flag_start3 <= '0'; 
   elsif pc_aux = "010101" then  
    flag_start2 <= '1'; 
    flag_start3 <= '0'; 
    flag_start1 <= '0'; 
   elsif pc_aux = "100001" then  
    flag_start3 <= '1'; 
    flag_start1 <= '0'; 
    flag_start2 <= '0'; 
   end if; 
  end if; 
 end process; 
  
 --Componentes 
 Comp1 : Memoria_Instrucciones port map( 
  input => pc_aux, 
  output => rom_output_aux 
 ); 
  
 Comp2 : Unidad_Ejecucion port map( 
  input_ex => rom_output_aux, 
  output_ex => output_ex_aux, 
  flag_zero => flag_zero_aux, 
  flag_signo => flag_signo_aux, 
  flag_acarreo => flag_acarreo_aux, 
  flag_overflow => flag_overflow_aux 
 ); 
  
 Comp3 : Converti port map( 
  S => "00" & output_ex_aux, 
  output_bcd => output_bcd_aux 
 ); 
  
 Comp4 : Parte2 port map( 
  input => output_bcd_aux(3 downto 0), 
  output => output_uni_aux 
 ); 
 
 Comp5 : Parte2 port map( 
  input => output_bcd_aux(7 downto 4), 
  output => output_dec_aux 
 ); 
 
 Comp6 : Parte2 port map( 
  input => output_bcd_aux(11 downto 8), 
  output => output_cen_aux 
 ); 
  
 Comp7 : Parte2 port map( 
  input => output_bcd_aux(15 downto 12), 
  output => output_mil_aux 
 ); 
  
 process(clk) 
 begin 
  if rising_edge(clk) then  
   if cuenta < 10000 then  
    cuenta <= cuenta + 1; 
   else 
    Seleccion <= Seleccion + 1; 
    cuenta <= 0; 
   end if; 
  end if; 
 end process; 
  
 --Mostrando displays 
 process(Seleccion) 
 begin 
  case Seleccion is 
   when "00" => 
    Mostrar <= "1110"; 
   when "01" => 
    Mostrar <= "1101"; 
   when "10" => 
    Mostrar <= "1011"; 
   when "11" =>  
    Mostrar <= "0111"; 
   when others =>  
    Mostrar <= "1111"; 
  end case; 
   
  case Mostrar is  
   when "1110" => 
    Segmentos <= output_uni_aux; 
   when "1101" => 
    Segmentos <= output_dec_aux; 
   when "1011" => 
    Segmentos <= output_cen_aux; 
   when "0111" =>  
    Segmentos <= output_mil_aux; 
   when others => 
    Segmentos <= "11111111"; 
end case; 
end process; 
Displays <= Mostrar; 
end architecture;