library ieee; 
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all; 
use ieee.numeric_std.all; 

entity Memoria_Instrucciones is 
    port( 
        input : in std_logic_vector(5 downto 0);
        output : out std_logic_vector(23 downto 0)
    );
end entity; 

architecture behavioral of Memoria_Instrucciones is
    
    -- ============================================
    -- MAPA DE OPCODES (SIN CONFLICTOS)
    -- ============================================
    -- PROGRAMA 1: 000000 - 001011
    -- PROGRAMA 2: 010000 - 011011  
    -- PROGRAMA 3: 100000 - 101011
    -- CONTROL:    111110 (WAIT_5S), 111111 (HALT)
    -- LECTURA:    110001, 110010, 110011
    -- ============================================
    
    type Rom_instrucciones is array(0 to 63) of std_logic_vector(23 downto 0);
    constant TR : Rom_instrucciones := ( 
        -- ====================================
        -- PROGRAMA 1: Direcciones 0-11
        -- Resultado: (13*X + 23*Y) * (W/4) = (39 + 138) * 2 = 354
        -- ====================================
        0  => "000000" & "000000" & "000000000000",  -- 13 * X → RAM[1]
        1  => "000001" & "000001" & "000000000000",  -- 23 * Y → RAM[2]
        2  => "000010" & "000010" & "000000000000",  -- W / 4  → RAM[3]
        3  => "000011" & "000011" & "000000000000",  -- Leer RAM[1] → dato1
        4  => "000100" & "000100" & "000000000000",  -- Leer RAM[2] → dato2
        5  => "000101" & "000101" & "000000000000",  -- dato1 + dato2 → RAM[1]
        6  => "000110" & "000110" & "000000000000",  -- Leer RAM[1] → dato1
        7  => "000111" & "000111" & "000000000000",  -- Leer RAM[3] → dato2
        8  => "001000" & "001000" & "000000000000",  -- dato1 * dato2 → RAM[1]
        9  => "110001" & "000000" & "000000000001",  -- LEER RESULTADO P1 (RAM[1])
        10 => "111110" & "000000" & "000000000000",  -- WAIT 5 SEGUNDOS
        11 => "111111" & "000000" & "000000000000",  -- HALT
        
        -- ====================================
        -- PROGRAMA 2: Direcciones 12-23
        -- Resultado: (X² * 13 + 30*X) - (Z/2) = (117 + 90) - 4 = 203
        -- ====================================
        12 => "010000" & "010000" & "000000000000",  -- X * X → RAM[1]
        13 => "010001" & "010001" & "000000000000",  -- Leer RAM[1] → dato1
        14 => "010010" & "010010" & "000000000000",  -- dato1 * 13 → RAM[1]
        15 => "010011" & "010011" & "000000000000",  -- 30 * X → RAM[2]
        16 => "010100" & "010100" & "000000000000",  -- Z / 2 → RAM[3]
        17 => "010101" & "010101" & "000000000000",  -- Leer RAM[1] → dato1
        18 => "010110" & "010110" & "000000000000",  -- Leer RAM[2] → dato2
        19 => "010111" & "010111" & "000000000000",  -- dato1 + dato2 → RAM[2]
        20 => "011000" & "011000" & "000000000000",  -- Leer RAM[2] → dato1
        21 => "011001" & "011001" & "000000000000",  -- Leer RAM[3] → dato2
        22 => "011010" & "011010" & "000000000000",  -- dato1 - dato2 → RAM[1]
        23 => "110010" & "000000" & "000000000001",  -- LEER RESULTADO P2 (RAM[1])
        24 => "111110" & "000000" & "000000000000",  -- WAIT 5 SEGUNDOS
        25 => "111111" & "000000" & "000000000000",  -- HALT
        
        -- ====================================
        -- PROGRAMA 3: Direcciones 26-37
        -- Resultado: (7*X² + 5*Z) - (W/5) = (63 + 40) - 2 = 101
        -- ====================================
        26 => "100000" & "100000" & "000000000000",  -- X * X → RAM[1]
        27 => "100001" & "100001" & "000000000000",  -- Leer RAM[1] → dato1
        28 => "100010" & "100010" & "000000000000",  -- dato1 * 7 → RAM[1]
        29 => "100011" & "100011" & "000000000000",  -- 5 * Z → RAM[2]
        30 => "100100" & "100100" & "000000000000",  -- W / 5 → RAM[3]
        31 => "100101" & "100101" & "000000000000",  -- Leer RAM[1] → dato1
        32 => "100110" & "100110" & "000000000000",  -- Leer RAM[2] → dato2
        33 => "100111" & "100111" & "000000000000",  -- dato1 + dato2 → RAM[2]
        34 => "101000" & "101000" & "000000000000",  -- Leer RAM[2] → dato1
        35 => "101001" & "101001" & "000000000000",  -- Leer RAM[3] → dato2
        36 => "101010" & "101010" & "000000000000",  -- dato1 - dato2 → RAM[3]
        37 => "110011" & "000000" & "000000000011",  -- LEER RESULTADO P3 (RAM[3])
        38 => "111110" & "000000" & "000000000000",  -- WAIT 5 SEGUNDOS
        39 => "111111" & "000000" & "000000000000",  -- HALT
        
        others => "111111" & "000000" & "000000000000"  -- HALT por defecto
    );
    
begin
    output <= TR(to_integer(unsigned(input))); 
end architecture;